library ieee;
     use ieee.std_logic_1164.all;

 entity up_counter is
     port (
         cout   :out integer := 0; -- Output of the counter
         enable :in  std_logic;                     -- Enable counting
         clk    :in  std_logic;                     -- Input clock
         reset  :in  std_logic                      -- Input reset
     );
 end entity;

architecture rtl of up_counter is
    signal coutTemp : integer := 0;
begin
     process (clk, reset) begin
         if (reset = '1') then
             coutTemp <= 0;
         elsif (rising_edge(clk)) then
             if (enable = '1') then
                 coutTemp <= coutTemp + 1;
             end if;
         end if;
         cout <= coutTemp;
     end process;
end architecture;
